module i_cache (
    input wire clk, rst,
    //mips core
    input         cpu_inst_req     ,
    input         cpu_inst_wr      ,
    input  [1 :0] cpu_inst_size    ,
    input  [31:0] cpu_inst_addr    ,
    input  [31:0] cpu_inst_wdata   ,
    output [31:0] cpu_inst_rdata   ,
    output        cpu_inst_addr_ok ,
    output        cpu_inst_data_ok ,

    //axi interface
    output         cache_inst_req     ,
    output         cache_inst_wr      ,
    output  [1 :0] cache_inst_size    ,
    output  [31:0] cache_inst_addr    ,
    output  [31:0] cache_inst_wdata   ,
    input   [31:0] cache_inst_rdata   ,
    input          cache_inst_addr_ok ,
    input          cache_inst_data_ok 
);
    //Cache配置
    parameter  INDEX_WIDTH  = 10, OFFSET_WIDTH = 2;
    localparam TAG_WIDTH    = 32 - INDEX_WIDTH - OFFSET_WIDTH;
    localparam CACHE_DEEPTH = 1 << INDEX_WIDTH;
    
    //Cache存储单元1
    reg                 cache_valid1 [CACHE_DEEPTH - 1 : 0];
    // reg                 cache_dirty1 [CACHE_DEEPTH - 1 : 0];
    reg [TAG_WIDTH-1:0] cache_tag1   [CACHE_DEEPTH - 1 : 0];
    reg [31:0]          cache_block1 [CACHE_DEEPTH - 1 : 0];

    //Cache存储单元2
    reg                 cache_valid2 [CACHE_DEEPTH - 1 : 0];
    // reg                 cache_dirty2 [CACHE_DEEPTH - 1 : 0];
    reg [TAG_WIDTH-1:0] cache_tag2   [CACHE_DEEPTH - 1 : 0];
    reg [31:0]          cache_block2 [CACHE_DEEPTH - 1 : 0];
    
    //访问地址分解
    wire [OFFSET_WIDTH-1:0] offset;
    wire [INDEX_WIDTH-1:0] index;
    wire [TAG_WIDTH-1:0] tag;
    
    assign offset = cpu_inst_addr[OFFSET_WIDTH - 1 : 0];
    assign index = cpu_inst_addr[INDEX_WIDTH + OFFSET_WIDTH - 1 : OFFSET_WIDTH];
    assign tag = cpu_inst_addr[31 : INDEX_WIDTH + OFFSET_WIDTH];

    //判断是否命中
    wire hit, hit1, hit2, miss;
    wire [31:0] c_block;
    assign hit1 = cache_valid1[index] & (cache_tag1[index] == tag);  //cache line1的valid位为1，且tag与地址中tag相等
    assign hit2 = cache_valid2[index] & (cache_tag2[index] == tag);  //cache line2的valid位为1，且tag与地址中tag相等
    assign hit = hit1 | hit2;
    assign miss = ~hit;
    assign c_block = hit1 ? cache_block1[index] : cache_block2[index];
    
    //FSM
    parameter IDLE = 2'b00, RM = 2'b01; // i cache只有read
    reg [1:0] state;
    always @(posedge clk) begin
        if(rst) begin
            state <= IDLE;
        end
        else begin
            case(state)
                IDLE:   state <= cpu_inst_req & miss ? RM : IDLE;
                RM:     state <= cache_inst_data_ok ? IDLE : RM;
            endcase
        end
    end

    //读内存
    //变量read_req, addr_rcv, read_finish用于构造类sram信号。
    wire read_req;      //一次完整的读事务，从发出读请求到结束
    reg addr_rcv;       //地址接收成功(addr_ok)后到结束
    wire read_finish;   //数据接收成功(data_ok)，即读请求结束
    always @(posedge clk) begin
        addr_rcv <= rst ? 1'b0 :
                    cache_inst_req & cache_inst_addr_ok ? 1'b1 :
                    read_finish ? 1'b0 : addr_rcv;
    end
    assign read_req = state==RM;
    assign read_finish = cache_inst_data_ok;

    //output to mips core
    assign cpu_inst_rdata   = hit ? c_block : cache_inst_rdata;
    assign cpu_inst_addr_ok = cpu_inst_req & hit | cache_inst_req & cache_inst_addr_ok;
    assign cpu_inst_data_ok = cpu_inst_req & hit | cache_inst_data_ok;

    //output to axi interface
    assign cache_inst_req   = read_req & ~addr_rcv;
    assign cache_inst_wr    = cpu_inst_wr;
    assign cache_inst_size  = cpu_inst_size;
    assign cache_inst_addr  = cpu_inst_addr;
    assign cache_inst_wdata = cpu_inst_wdata;

    //写入Cache
    //保存地址中的tag, index，防止addr发生改变
    reg [TAG_WIDTH-1:0] tag_save;
    reg [INDEX_WIDTH-1:0] index_save;
    reg group_save;
    always @(posedge clk) begin
        tag_save   <= rst ? 0 :
                      cpu_inst_req ? tag : tag_save;
        index_save <= rst ? 0 :
                      cpu_inst_req ? index : index_save;
        group_save <= rst ? 0 :
                      cpu_inst_req ? ((~cache_valid1[index] || cache_valid2[index]) ? 1'b0 : 1'b1) : group_save;
    end

    integer t;
    always @(posedge clk) begin
        if(rst) begin
            for(t=0; t<CACHE_DEEPTH; t=t+1) begin   //刚开始将Cache置为无效
                cache_valid1[t] <= 0;
                cache_valid2[t] <= 0;
            end
        end
        else begin
            if(read_finish) begin //读缺失，访存结束时
                if(group_save) begin    
                    cache_valid2[index_save] <= 1'b1;             //将Cache line置为有效
                    cache_tag2  [index_save] <= tag_save;
                    cache_block2[index_save] <= cache_inst_rdata; //写入Cache line
                end
                else begin
                    cache_valid1[index_save] <= 1'b1;             //将Cache line置为有效
                    cache_tag1  [index_save] <= tag_save;
                    cache_block1[index_save] <= cache_inst_rdata; //写入Cache line
                end
            end
        end
    end
endmodule